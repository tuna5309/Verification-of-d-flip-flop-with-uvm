class d_sequencer extends uvm_sequencer#(df_data);
	`uvm_component_utils(d_sequencer)
	
	function new (string name = "d_sequencer ",uvm_component parent);
		super.new(name);
	endfunction
	
	
	

endclass 
