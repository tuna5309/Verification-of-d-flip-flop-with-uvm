interface df_intf;
	logic clk,reset;
	logic d;
	logic q_out;
endinterface 


